** Profile: "SCHEMATIC1-Q_point"  [ C:\Users\EMTOO\Desktop\Papers\p1-schematic1-q_point.sim ] 

** Creating circuit file "p1-schematic1-q_point.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 1 1000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "..\..\..\public\music\p1-SCHEMATIC1.net" 


.END
