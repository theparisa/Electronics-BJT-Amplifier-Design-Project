** Profile: "SCHEMATIC1-p4_sim"  [ C:\Users\Public\Music\p4-SCHEMATIC1-p4_sim.sim ] 

** Creating circuit file "p4-SCHEMATIC1-p4_sim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB ".\p4.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 10 10k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p4-SCHEMATIC1.net" 


.END
