** Profile: "SCHEMATIC1-sim_3"  [ C:\Users\Public\Music\p3-SCHEMATIC1-sim_3.sim ] 

** Creating circuit file "p3-SCHEMATIC1-sim_3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10 10 10k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\p3-SCHEMATIC1.net" 


.END
